module AND_GATE
(
input A, B,
output C
);
assign C = A&B;
endmodule 